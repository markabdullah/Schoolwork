module vga

end module
